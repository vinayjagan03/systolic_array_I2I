`ifndef SYSTOLIC_ARRAY_PKG_SVH
`define SYSTOLIC_ARRAY_PKG_SVH

localparam WORD_SIZE = 32;

typedef logic [WORD_SIZE-1:0] word_t;

`endif // SYSTOLIC_ARRAY_PKG_SVH