module top_systolic_array (
    input logic clk, n_rst,
    input logic start_matmul,
    output logic done
);


    
endmodule