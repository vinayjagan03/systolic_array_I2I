module fp32 (
    input logic clk, n_rst,
    input word_t a,
    input word_t b,
    input word_t c,
    input logic start_mac,
    output logic ready,
    output word_t result
);
    
endmodule