`include "systolic_array_pkg.svh"

module fp32_stage_mantissa_mul (
    input logic clk, n_rst,
    input logic valid_i,
    input logic [22:0] mantissa_a,
    input logic [22:0] mantissa_b,
    input logic [9:0] exponent_sum,
    input logic sign,

);
    
endmodule